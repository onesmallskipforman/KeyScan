module shiftreg #(parameter N = 8)
					  (input logic clk,
						input logic reset, load,
						input logic sin)